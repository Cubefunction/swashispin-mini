`timescale 1ns / 1ps

module uart_api_dc
#(parameter DAC_WIDTH=16,
     parameter CYCLE_WIDTH=30,
     parameter DAC_CHANNEL=24,
     parameter CHANNEL_MES_WIDTH=96,
     parameter STREAM_ITER_WIDTH=10,
     parameter CORE_ITER_WIDTH=10,
     parameter DEPTH=10,
     parameter INSN_WIDTH=DAC_WIDTH*2+CORE_ITER_WIDTH+CYCLE_WIDTH,
     parameter TOTAL_REGS=DEPTH*3+2)
     (input  logic i_clk, i_rst,

     input  logic i_rx,
     output logic o_tx,

     //input  logic i_trigger,
     
     output logic [DAC_CHANNEL-1:0] o_sclk,
     output logic [DAC_CHANNEL-1:0]o_mosi,
     output logic [DAC_CHANNEL-1:0]o_cs_n,
     output logic [DAC_CHANNEL-1:0] o_ldac_n);

    logic w_deq_rxq, w_rxq_empty;
    logic [7:0] w_rxq_data;
    
    localparam NUM_BYTES = INSN_WIDTH / 8;
    localparam FRAME_BYTES = 62 * 4; 
    localparam FRAME_WORDS = 62;
    
    uart #(
        .DATA_WIDTH(8),
        .RX_FIFO_DEPTH(100),
        .RX_FIFO_AF_DEPTH(16),
        .RX_FIFO_AE_DEPTH(4),
        .TX_FIFO_DEPTH(20),
        .TX_FIFO_AF_DEPTH(16),
        .TX_FIFO_AE_DEPTH(4)
    ) U (
        .i_clk(i_clk),
        .i_rst(!i_rst),
        .i_rx(i_rx),
        .o_tx(o_tx),
        .i_deq_rxq(w_deq_rxq),
        .o_rxq_data(w_rxq_data),
        .o_rxq_empty(w_rxq_empty),
        /* verilator lint_off PINCONNECTEMPTY */
        .o_rxq_ae(),
        .o_rxq_full(),
        .o_rxq_af(),
        .i_enq_txq(),
        .i_txq_data(),
        .o_txq_empty(),
        .o_txq_ae(),
        .o_txq_full(),
        .o_txq_af()
    );

    assign w_deq_rxq = !w_rxq_empty;
// ================================================================
// UART-----FIFO32 
// ================================================================
    logic [1:0]  r_byte_cnt;
    logic [31:0] r_word_buf;
    logic        w_fifo32_enq;

     always_ff @(posedge i_clk or negedge i_rst) begin
        if (!i_rst) begin
            r_byte_cnt   <= 'd0;
            r_word_buf   <= 'd0;
            w_fifo32_enq <= 1'b0;
        end
        else if (!w_rxq_empty) begin
            r_word_buf <= {r_word_buf[23:0],w_rxq_data };
    
            if (r_byte_cnt == 'd3) begin
                w_fifo32_enq <= 1'b1;   // write FIFO32
                r_byte_cnt   <= 'd0;
            end
            else begin
                w_fifo32_enq <= 1'b0;
                r_byte_cnt   <= r_byte_cnt + 'd1;
            end
        end
        else begin
            w_fifo32_enq <= 1'b0;  
        end
    end

// ================================================================
// 32-bit FIFO 
// ================================================================

    logic        w_fifo32_full, w_fifo32_empty;
    logic [31:0] w_fifo32_dout;
    logic        w_fifo32_deq;

    fifo #(
        .WIDTH(32),
        .DEPTH(64),       
        .AF_DEPTH(56),
        .AE_DEPTH(8)
    ) u_fifo32 (
        .i_clk(i_clk),
        .i_rst(!i_rst),
        .i_data(r_word_buf),
        .i_enq(w_fifo32_enq),
        .i_deq(w_fifo32_deq),   
        .o_data(w_fifo32_dout),
        .o_full(w_fifo32_full),
        .o_empty(w_fifo32_empty),
        .o_almost_full(),
        .o_almost_empty()
    );
// ================================================================
// 62*32 register from fifo
// ================================================================

    dc_dispatcher #(
        .DAC_CHANNEL(DAC_CHANNEL),
        .FRAME_WORDS(TOTAL_REGS)
    ) u_dispatcher (
        .i_clk(i_clk),
        .i_rst(i_rst),
        .i_fifo_data(w_fifo32_dout),
        .i_fifo_empty(w_fifo32_empty),
        .o_fifo_deq(w_fifo32_deq),
        .o_dc_regs(w_dc_regs),
        .o_channel_sel(w_channel_sel),
        .o_valid_frame(w_valid_frame),
        .o_launch_cmd(w_launch_cmd_reg)
    );

    logic [61:0][31:0]   w_dc_regs;       
    logic [4:0]          w_channel_sel;   
    logic                w_valid_frame; 
    logic [3:0][31:0]    w_launch_cmd_reg;

    logic [DAC_CHANNEL-1:0][61:0][31:0] r_dc_regs;  
    logic [DAC_CHANNEL-1:0]             r_start;     
    logic [DAC_CHANNEL-1:0]             w_armed;     


    always_ff @(posedge i_clk or negedge i_rst) begin
    if (!i_rst) begin
        r_dc_regs <= '0;
    end else if (w_valid_frame) begin
        case (w_channel_sel)
            5'd0 :  r_dc_regs[0]  <= w_dc_regs;
            5'd1 :  r_dc_regs[1]  <= w_dc_regs;
            5'd2 :  r_dc_regs[2]  <= w_dc_regs;
            5'd3 :  r_dc_regs[3]  <= w_dc_regs;
            5'd4 :  r_dc_regs[4]  <= w_dc_regs;
            5'd5 :  r_dc_regs[5]  <= w_dc_regs;
            5'd6 :  r_dc_regs[6]  <= w_dc_regs;
            5'd7 :  r_dc_regs[7]  <= w_dc_regs;
            5'd8 :  r_dc_regs[8]  <= w_dc_regs;
            5'd9 :  r_dc_regs[9]  <= w_dc_regs;
            5'd10:  r_dc_regs[10] <= w_dc_regs;
            5'd11:  r_dc_regs[11] <= w_dc_regs;
            5'd12:  r_dc_regs[12] <= w_dc_regs;
            5'd13:  r_dc_regs[13] <= w_dc_regs;
            5'd14:  r_dc_regs[14] <= w_dc_regs;
            5'd15:  r_dc_regs[15] <= w_dc_regs;
            5'd16:  r_dc_regs[16] <= w_dc_regs;
            5'd17:  r_dc_regs[17] <= w_dc_regs;
            5'd18:  r_dc_regs[18] <= w_dc_regs;
            5'd19:  r_dc_regs[19] <= w_dc_regs;
            5'd20:  r_dc_regs[20] <= w_dc_regs;
            5'd21:  r_dc_regs[21] <= w_dc_regs;
            5'd22:  r_dc_regs[22] <= w_dc_regs;
            5'd23:  r_dc_regs[23] <= w_dc_regs;
            default: ;
        endcase
    end
end
   genvar i;
   generate
       for (i = 0; i < DAC_CHANNEL; i++) begin : GEN_DC
           dc #(
               .DAC_WIDTH(DAC_WIDTH),
               .CYCLE_WIDTH(CYCLE_WIDTH),
               .STREAM_ITER_WIDTH(STREAM_ITER_WIDTH),
               .CORE_ITER_WIDTH(CORE_ITER_WIDTH),
               .DEPTH(DEPTH)
           ) u_dc (
               .i_clk(i_clk),
               .i_rst(i_rst),
               .i_regs(r_dc_regs[i]),
               .i_start(r_start[i]),
               .o_armed(w_armed[i]),
               .o_sclk(o_sclk[i]),
               .o_mosi(o_mosi[i]),
               .o_cs_n(o_cs_n[i]),
               .o_ldac_n(o_ldac_n[i])
           );
       end
   endgenerate

    
   launch #(
    .NUM_DC_CHANNEL(24),
    .NUM_RF_CHANNEL(7),
    .NUM_LI_CHANNEL(2)
    )u_launch(
       .i_clk(i_clk), 
       .i_rst(i_rst),

       .i_regs(w_launch_cmd_reg),

       .i_dc_armed(w_armed),
       //.i_rf_armed(),
       //.i_li_armed(),

       .o_dc_start(r_start)
       //.o_rf_start(),
       //.o_li_start()
       );



endmodule
